grammar edu:umn:cs:melt:exts:ableC:attributeGrammars:concretesyntax;

imports edu:umn:cs:melt:ableC:concretesyntax;
imports silver:langutil only ast; 

imports edu:umn:cs:melt:exts:ableC:attributeGrammars:abstractsyntax;
