grammar edu:umn:cs:melt:exts:ableC:attributeGrammars:abstractsyntax;

